library verilog;
use verilog.vl_types.all;
entity Ripple_Adder_4bit_vlg_vec_tst is
end Ripple_Adder_4bit_vlg_vec_tst;
