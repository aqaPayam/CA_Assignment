library verilog;
use verilog.vl_types.all;
entity Adder64Bit_vlg_vec_tst is
end Adder64Bit_vlg_vec_tst;
