library verilog;
use verilog.vl_types.all;
entity FinalCircuit_vlg_vec_tst is
end FinalCircuit_vlg_vec_tst;
