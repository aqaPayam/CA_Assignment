library verilog;
use verilog.vl_types.all;
entity BarrelShifter8Bit_vlg_vec_tst is
end BarrelShifter8Bit_vlg_vec_tst;
