library verilog;
use verilog.vl_types.all;
entity Adder32BIt_vlg_vec_tst is
end Adder32BIt_vlg_vec_tst;
