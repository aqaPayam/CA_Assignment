library verilog;
use verilog.vl_types.all;
entity Adder12Bit_vlg_vec_tst is
end Adder12Bit_vlg_vec_tst;
