library verilog;
use verilog.vl_types.all;
entity CarrySelectAdder16Bit_vlg_vec_tst is
end CarrySelectAdder16Bit_vlg_vec_tst;
