library verilog;
use verilog.vl_types.all;
entity Multiplier4Bits_vlg_vec_tst is
end Multiplier4Bits_vlg_vec_tst;
