library verilog;
use verilog.vl_types.all;
entity CarrySkipAdder4Bit_vlg_vec_tst is
end CarrySkipAdder4Bit_vlg_vec_tst;
