library verilog;
use verilog.vl_types.all;
entity CarrySkipAdder16Bit_vlg_vec_tst is
end CarrySkipAdder16Bit_vlg_vec_tst;
