library verilog;
use verilog.vl_types.all;
entity ClaFourBitAdder_vlg_vec_tst is
end ClaFourBitAdder_vlg_vec_tst;
