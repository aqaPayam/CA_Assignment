library verilog;
use verilog.vl_types.all;
entity BusMux_vlg_vec_tst is
end BusMux_vlg_vec_tst;
